typedef class environment;
event clock_env , reset_env;

//interface testSignals();
interface testSignals(input clock, input resetb);
  logic test1;
endinterface
