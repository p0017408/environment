`include "interface.sv"
`include "clkrst_monitor.sv"
`include "seqer.sv"
`include "bfm.sv"
